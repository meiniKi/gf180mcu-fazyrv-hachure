VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_hachure_ip__logo
  CLASS BLOCK ;
  FOREIGN gf180mcu_hachure_ip__logo ;
  ORIGIN 0.000 0.000 ;
  SIZE 225 BY 375 ;
  OBS
      LAYER Metal5 ;
        RECT 0.0 0.0 225 375 ;
  END
END gf180mcu_hachure_ip__logo
END LIBRARY

