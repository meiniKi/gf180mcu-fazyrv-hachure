module gf180mcu_fazyrv_ip__logo;
endmodule
