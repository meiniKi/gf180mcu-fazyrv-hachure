module gf180mcu_hachure_ip__logo;
endmodule
